module control (
    //main decoder
    input logic [6:0] op_code,
    input logic zero,
    output logic [2:0] imm_type,
    output logic mem_write,
    output logic reg_write,
    output logic alu_source,
    output logic result_source,

    //alu decoder
    input  logic [2:0] func3,
    input  logic [6:0] func7,
    output logic [2:0] alu_control
);


  logic [1:0] alu_op;

  always_comb begin : MAIN_DECODER
    case (op_code)
      // I-type
      7'b0000011: begin
        imm_type = 3'b000;
        mem_write = 1'b0;
        reg_write = 1'b1;
        alu_op = 2'b00;
        alu_source = 1'b1;
        result_source = 1'b1;
      end

      // S-type
      7'b0100011: begin
        imm_type = 3'b001;
        mem_write = 1'b1;
        reg_write = 1'b0;
        alu_op = 2'b00;
        alu_source = 1'b1;
      end

      //R-type
      7'b0110011: begin
        mem_write = 1'b0;
        reg_write = 1'b1;
        alu_op = 2'b10;
        alu_source = 1'b0;
        result_source = 1'b0;
      end

      default: begin
        imm_type = 3'b000;
        mem_write = 1'b0;
        reg_write = 1'b0;
        alu_op = 2'b11;
      end
    endcase
  end


  always_comb begin : ALU_DECODER
    case (alu_op)
      // LW, SW
      2'b00:   alu_control = 3'b000;
      // R-type
      2'b10: begin
        case (func3)
          // ADD
          3'b000: alu_control = 3'b000;
          // OR
          3'b110: alu_control = 3'b011;
          // AND
          3'b111: alu_control = 3'b010;

          default: alu_control = 3'b111;
        endcase
      end
      default: alu_control = 3'b111;
    endcase
  end

endmodule
